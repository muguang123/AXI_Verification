package axi_test_pkg;

	import uvm_pkg::*;
	
	`include "uvm_macros.svh"
	`include "master_xtn.sv"
	`include "master_agt_cfg.sv"
	`include "slave_agt_cfg.sv"
	`include "axi_env_config.sv"
	`include "master_driver.sv"
	`include "master_sequencer.sv"
	`include "master_monitor.sv"
	`include "master_agent.sv"
	`include "master_agt_top.sv"
	`include "master_sequence.sv"
	`include "slave_xtn.sv"
	`include "slave_sequencer.sv"
	`include "slave_monitor.sv"
	`include "slave_sequence.sv"
	`include "slave_driver.sv"
	`include "slave_agent.sv"
	`include "slave_agt_top.sv"
	`include "virtual_sequencer.sv"
	`include "axi_virtual_seq.sv"
	`include "axi_scoreboard.sv"
	`include "avi_environment.sv"
	`include "axi_test.sv"


endpackage
